package shared_pkg;
    int test_finished;
    int error_count_out = 0, correct_count_out = 0;
    int error_count_ack = 0, correct_count_ack = 0;
    int error_count_over = 0, correct_count_over = 0;
    int error_count_full = 0, correct_count_full = 0;
    int error_count_empty = 0, correct_count_empty = 0;
    int error_count_almostfull = 0, correct_count_almostfull = 0;
    int error_count_almostempty = 0, correct_count_almostempty = 0;
    int error_count_under = 0, correct_count_under = 0;
endpackage